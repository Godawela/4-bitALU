<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-82.619,26.904,246.422,-138.796</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>16.5,-15.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>16.5,-20</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>37,-16</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>27,-20</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AO_XNOR2</type>
<position>56.5,-13</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>37,-24</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_SMALL_INVERTER</type>
<position>27,-23</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>73.5,-14</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND3</type>
<position>73.5,-26.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_OR4</type>
<position>92.5,-11.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>38 </input>
<input>
<ID>IN_3</ID>39 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>12,-39</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>12,-48</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>34,-37.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>34,-47</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,-41</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_SMALL_INVERTER</type>
<position>24.5,-44.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AO_XNOR2</type>
<position>48,-41.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>10,-60</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>10,-75.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>28,-61</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>28.5,-75</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_SMALL_INVERTER</type>
<position>19,-67.5</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_SMALL_INVERTER</type>
<position>19.5,-72.5</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AO_XNOR2</type>
<position>44,-64</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND4</type>
<position>84.5,-55.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>26 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>9,-88.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>9.5,-100</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>27.5,-89.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND2</type>
<position>27.5,-99</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AE_SMALL_INVERTER</type>
<position>17.5,-93</position>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_SMALL_INVERTER</type>
<position>18.5,-96.5</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AO_XNOR2</type>
<position>42.5,-94.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>93.5,-84.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND3</type>
<position>88,-104.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>20 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND4</type>
<position>88.5,-144</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>28 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_OR4</type>
<position>112.5,-88.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>40 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>34 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND4</type>
<position>80,-112.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>24 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>103,-11</position>
<input>
<ID>N_in0</ID>41 </input>
<input>
<ID>N_in1</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>121,-88</position>
<input>
<ID>N_in0</ID>42 </input>
<input>
<ID>N_in2</ID>42 </input>
<input>
<ID>N_in3</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>99.5,-144</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>10,-14.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>10,-19</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>5.5,-38</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>5,-46.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>4.5,-60.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>4,-75</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>3.5,-88</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>3.5,-99</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>107,-8.5</position>
<gparam>LABEL_TEXT L</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>126.5,-87</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>105.5,-143.5</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-15.5,31,-15.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>23.5 4</intersection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-15.5,31,-4</points>
<intersection>-15.5 1</intersection>
<intersection>-15 8</intersection>
<intersection>-4 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>23.5,-23,23.5,-15.5</points>
<intersection>-23 5</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>23.5,-23,25,-23</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>23.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>31,-4,87,-4</points>
<intersection>31 3</intersection>
<intersection>87 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>87,-8.5,87,-4</points>
<intersection>-8.5 9</intersection>
<intersection>-4 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>31,-15,34,-15</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>31 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>87,-8.5,89.5,-8.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>87 7</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-20,25,-20</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>22 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>22,-25,22,-20</points>
<intersection>-25 6</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>22,-25,34,-25</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>22 5</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-20,31.5,-17</points>
<intersection>-20 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-17,34,-17</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-20,31.5,-20</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-16,46.5,-12</points>
<intersection>-16 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-12,53.5,-12</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-16,46.5,-16</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-23,34,-23</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-34,50,-14</points>
<intersection>-34 3</intersection>
<intersection>-24 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-14,53.5,-14</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-24,50,-24</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50,-34,105.5,-34</points>
<intersection>50 0</intersection>
<intersection>105.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>105.5,-85.5,105.5,-34</points>
<intersection>-85.5 5</intersection>
<intersection>-34 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>105.5,-85.5,109.5,-85.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>105.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-13,70.5,-13</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-141,67,-13</points>
<intersection>-141 13</intersection>
<intersection>-102.5 11</intersection>
<intersection>-83.5 9</intersection>
<intersection>-52.5 6</intersection>
<intersection>-24.5 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67,-24.5,70.5,-24.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>67,-52.5,81.5,-52.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>67,-83.5,90.5,-83.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>67,-102.5,85,-102.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection>
<intersection>75.5 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>67,-141,85.5,-141</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>67 3</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>75.5,-109.5,75.5,-102.5</points>
<intersection>-109.5 15</intersection>
<intersection>-102.5 11</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>75.5,-109.5,77,-109.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>75.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-44.5,18,-36.5</points>
<intersection>-44.5 3</intersection>
<intersection>-39 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-36.5,31,-36.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-39,18,-39</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>18,-44.5,22.5,-44.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-48,31,-48</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>19.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>19.5,-48,19.5,-41</points>
<intersection>-48 1</intersection>
<intersection>-41 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>19.5,-41,24,-41</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>19.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-41,28.5,-38.5</points>
<intersection>-41 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-38.5,31,-38.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-41,28.5,-41</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-46,28.5,-44.5</points>
<intersection>-46 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-46,31,-46</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-44.5,28.5,-44.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-37.5,62.5,-37.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>45 5</intersection>
<intersection>62.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62.5,-37.5,62.5,-15</points>
<intersection>-37.5 1</intersection>
<intersection>-15 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62.5,-15,70.5,-15</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>62.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>45,-40.5,45,-37.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-85.5,39,-42.5</points>
<intersection>-85.5 3</intersection>
<intersection>-47 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-42.5,45,-42.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-47,39,-47</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39,-85.5,90.5,-85.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-143,60.5,-26.5</points>
<intersection>-143 7</intersection>
<intersection>-104.5 5</intersection>
<intersection>-54.5 3</intersection>
<intersection>-41.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-26.5,70.5,-26.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-41.5,60.5,-41.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60.5,-54.5,81.5,-54.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>60.5,-104.5,85,-104.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection>
<intersection>71.5 8</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>60.5,-143,85.5,-143</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>71.5,-111.5,71.5,-104.5</points>
<intersection>-111.5 10</intersection>
<intersection>-104.5 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>71.5,-111.5,77,-111.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>71.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-60,25,-60</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-72.5,16,-60</points>
<intersection>-72.5 4</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,-72.5,17.5,-72.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-79,14.5,-67.5</points>
<intersection>-79 3</intersection>
<intersection>-75.5 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-67.5,17,-67.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-75.5,14.5,-75.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14.5,-79,23.5,-79</points>
<intersection>14.5 0</intersection>
<intersection>23.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>23.5,-79,23.5,-76</points>
<intersection>-79 3</intersection>
<intersection>-76 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>23.5,-76,25.5,-76</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>23.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-67.5,23,-62</points>
<intersection>-67.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-62,25,-62</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-67.5,23,-67.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-74,23.5,-72.5</points>
<intersection>-74 1</intersection>
<intersection>-72.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-74,25.5,-74</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-72.5,23.5,-72.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-61,70.5,-61</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>40 4</intersection>
<intersection>70.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-61,70.5,-28.5</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>40,-63,40,-61</points>
<intersection>-63 5</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>40,-63,41,-63</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>40 4</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-106.5,33,-65</points>
<intersection>-106.5 3</intersection>
<intersection>-75 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-65,41,-65</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-75,33,-75</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-106.5,85,-106.5</points>
<connection>
<GID>72</GID>
<name>IN_2</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-145,56.5,-56.5</points>
<intersection>-145 3</intersection>
<intersection>-113.5 4</intersection>
<intersection>-64 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-56.5,81.5,-56.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-64,56.5,-64</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>56.5,-145,85.5,-145</points>
<connection>
<GID>74</GID>
<name>IN_2</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>56.5,-113.5,77,-113.5</points>
<connection>
<GID>82</GID>
<name>IN_2</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-88.5,24.5,-88.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>14.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-96.5,14.5,-88.5</points>
<intersection>-96.5 4</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-96.5,16.5,-96.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-100,13.5,-93</points>
<intersection>-100 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-93,15.5,-93</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-100,24.5,-100</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-93,22,-90.5</points>
<intersection>-93 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-90.5,24.5,-90.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection>
<intersection>23.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-93,22,-93</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,-115.5,23.5,-90.5</points>
<intersection>-115.5 4</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23.5,-115.5,77,-115.5</points>
<connection>
<GID>82</GID>
<name>IN_3</name></connection>
<intersection>23.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-98,22.5,-96.5</points>
<intersection>-98 1</intersection>
<intersection>-96.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-98,24.5,-98</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-96.5,22.5,-96.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-89.5,75.5,-89.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>37 4</intersection>
<intersection>75.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-89.5,75.5,-58.5</points>
<intersection>-89.5 1</intersection>
<intersection>-58.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>37,-93.5,37,-89.5</points>
<intersection>-93.5 6</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>75.5,-58.5,81.5,-58.5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>75.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>37,-93.5,39.5,-93.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>37 4</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-99,35,-95.5</points>
<intersection>-99 2</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-95.5,39.5,-95.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-99,35,-99</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-147,49.5,-94.5</points>
<intersection>-147 1</intersection>
<intersection>-94.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-147,85.5,-147</points>
<connection>
<GID>74</GID>
<name>IN_3</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-94.5,49.5,-94.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-104.5,100,-91.5</points>
<intersection>-104.5 2</intersection>
<intersection>-91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-91.5,109.5,-91.5</points>
<connection>
<GID>80</GID>
<name>IN_3</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-104.5,100,-104.5</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-89.5,103,-84.5</points>
<intersection>-89.5 1</intersection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-89.5,109.5,-89.5</points>
<connection>
<GID>80</GID>
<name>IN_2</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-84.5,103,-84.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-14,82,-10.5</points>
<intersection>-14 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-10.5,89.5,-10.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-14,82,-14</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-26.5,83,-12.5</points>
<intersection>-26.5 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-12.5,89.5,-12.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-26.5,83,-26.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-55.5,88.5,-14.5</points>
<intersection>-55.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-14.5,89.5,-14.5</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-55.5,88.5,-55.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-112.5,96,-87.5</points>
<intersection>-112.5 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-112.5,96,-112.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96,-87.5,109.5,-87.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-11.5,104,-11.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>102 4</intersection>
<intersection>104 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>102,-11.5,102,-11</points>
<connection>
<GID>84</GID>
<name>N_in0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>104,-11.5,104,-11</points>
<connection>
<GID>84</GID>
<name>N_in1</name></connection>
<intersection>-11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-88.5,120,-88.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>120 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>120,-88.5,120,-87</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<intersection>-88.5 1</intersection>
<intersection>-87 8</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>121.5,-89,121.5,-87</points>
<intersection>-89 7</intersection>
<intersection>-87 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>121,-89,121.5,-89</points>
<connection>
<GID>86</GID>
<name>N_in2</name></connection>
<intersection>121.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>120,-87,121.5,-87</points>
<connection>
<GID>86</GID>
<name>N_in3</name></connection>
<intersection>120 3</intersection>
<intersection>121.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-144,98.5,-144</points>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 1>
<page 2>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 2>
<page 3>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 3>
<page 4>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 4>
<page 5>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 5>
<page 6>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 6>
<page 7>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 7>
<page 8>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 8>
<page 9>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 9></circuit>