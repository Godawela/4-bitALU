<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>5.24199,-8.72672,252.023,-133.002</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>45.5,-6.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-9.5,-111.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>58,-88.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>58,-101</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>58,-109.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>58.5,-71.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>59.5,-24.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_XOR2</type>
<position>72.5,-88</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AE_OR2</type>
<position>66,-104</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>76.5,-83.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>88.5,-6</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AI_XOR2</type>
<position>101.5,-88.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AI_XOR2</type>
<position>114,-88.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>101.5,-101</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>101.5,-109.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR2</type>
<position>115.5,-105</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AI_XOR2</type>
<position>102,-71.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>103,-23</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>118,-84</position>
<input>
<ID>N_in2</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>133.5,-3.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR2</type>
<position>146,-88</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AI_XOR2</type>
<position>158.5,-88</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>146,-100.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>146,-109</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_OR2</type>
<position>160,-104.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>146.5,-71</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>147.5,-20</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>162.5,-83.5</position>
<input>
<ID>N_in2</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>165.5,-104.5</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>-1,-7</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AI_XOR2</type>
<position>11.5,-93.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AI_XOR2</type>
<position>24,-93.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_AND2</type>
<position>11.5,-106</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>165.5,-107.5</position>
<gparam>LABEL_TEXT C3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>11.5,-114.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>118.5,-108.5</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AE_OR2</type>
<position>25.5,-110</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>69.5,-107.5</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AI_XOR2</type>
<position>12,-76.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>29.5,-112.5</position>
<gparam>LABEL_TEXT C0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>15.5,-20.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>-7,-7.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>28,-89</position>
<input>
<ID>N_in2</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>11,-20.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>104,-128.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>29 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>40.5,-6.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>56,-23.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>84,-6.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>99,-24</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>128.5,-5.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>142.5,-20</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>-13,-111</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>-12,-114.5</position>
<gparam>LABEL_TEXT Add 0 / Sub 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>28,-86</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>76,-81</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>115.5,-83.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>162,-81</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>206,-28.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_SMALL_INVERTER</type>
<position>196,-32.5</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AO_XNOR2</type>
<position>225.5,-25.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>206,-36.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_SMALL_INVERTER</type>
<position>196,-35.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>241,-25.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND3</type>
<position>242.5,-39</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_OR4</type>
<position>261.5,-24</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND2</type>
<position>203,-50</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_AND2</type>
<position>203,-59.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_SMALL_INVERTER</type>
<position>195,-53.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_SMALL_INVERTER</type>
<position>193.5,-57</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AO_XNOR2</type>
<position>217,-54</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_AND2</type>
<position>197,-73.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>197.5,-87.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_SMALL_INVERTER</type>
<position>188,-80</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_SMALL_INVERTER</type>
<position>188.5,-85</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AO_XNOR2</type>
<position>213,-76.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND4</type>
<position>253.5,-68</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>63 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND2</type>
<position>196.5,-102</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_AND2</type>
<position>196.5,-111.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_SMALL_INVERTER</type>
<position>186.5,-105.5</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AE_SMALL_INVERTER</type>
<position>187.5,-109</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>93</ID>
<type>AO_XNOR2</type>
<position>211.5,-107</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND2</type>
<position>262.5,-97</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND3</type>
<position>256.5,-117.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>57 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND4</type>
<position>257.5,-156.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>65 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_OR4</type>
<position>281.5,-101</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>67 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND4</type>
<position>249,-125</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>99</ID>
<type>GA_LED</type>
<position>272,-23.5</position>
<input>
<ID>N_in1</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>290,-100.5</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>GA_LED</type>
<position>268.5,-156.5</position>
<input>
<ID>N_in0</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>276,-21</position>
<gparam>LABEL_TEXT L</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>295.5,-99.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>274.5,-156</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-68.5,59.5,-26.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-62.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>59.5,-62.5,183,-62.5</points>
<intersection>59.5 0</intersection>
<intersection>183 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>183,-88.5,183,-62.5</points>
<intersection>-88.5 13</intersection>
<intersection>-80 14</intersection>
<intersection>-62.5 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>183,-88.5,194.5,-88.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>183 12</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>183,-80,186,-80</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>183 12</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-108.5,53.5,-76.5</points>
<intersection>-108.5 5</intersection>
<intersection>-87.5 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-87.5,55,-87.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-76.5,58.5,-76.5</points>
<intersection>53.5 0</intersection>
<intersection>58.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58.5,-76.5,58.5,-74.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>53.5,-108.5,55,-108.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-122.5,45.5,-8.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-122.5,82.5,-122.5</points>
<intersection>45.5 0</intersection>
<intersection>51 3</intersection>
<intersection>55 9</intersection>
<intersection>82.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,-122.5,51,-89.5</points>
<intersection>-122.5 1</intersection>
<intersection>-89.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>51,-89.5,55,-89.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>82.5,-136.5,82.5,-122.5</points>
<intersection>-136.5 10</intersection>
<intersection>-122.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>55,-122.5,55,-110.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>82.5,-136.5,174,-136.5</points>
<intersection>82.5 8</intersection>
<intersection>95.5 14</intersection>
<intersection>174 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>174,-136.5,174,-72.5</points>
<intersection>-136.5 10</intersection>
<intersection>-85 16</intersection>
<intersection>-72.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>174,-72.5,194,-72.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>174 12</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>95.5,-136.5,95.5,-128.5</points>
<intersection>-136.5 10</intersection>
<intersection>-128.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>95.5,-128.5,101,-128.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>95.5 14</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>174,-85,186.5,-85</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>174 12</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-93,64,-87</points>
<intersection>-93 2</intersection>
<intersection>-88.5 5</intersection>
<intersection>-87 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-93,64,-93</points>
<intersection>48.5 3</intersection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-102,48.5,-93</points>
<intersection>-102 7</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>61,-88.5,64,-88.5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>48.5,-102,55,-102</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>48.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>64,-87,69.5,-87</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-110,41.5,-96.5</points>
<intersection>-110 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-96.5,69.5,-96.5</points>
<intersection>41.5 0</intersection>
<intersection>52 4</intersection>
<intersection>69.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-110,41.5,-110</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69.5,-96.5,69.5,-89</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>52,-100,52,-96.5</points>
<intersection>-100 5</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>52,-100,55,-100</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>52 4</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-103,62,-101</points>
<intersection>-103 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-103,63,-103</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-101,62,-101</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-109.5,62,-105</points>
<intersection>-109.5 2</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-105,63,-105</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-109.5,62,-109.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-88,76,-83.5</points>
<intersection>-88 2</intersection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-83.5,76,-83.5</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-88,76,-88</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-104,108.5,-101</points>
<intersection>-104 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-104,112.5,-104</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-101,108.5,-101</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-109.5,108,-106</points>
<intersection>-109.5 2</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-106,112.5,-106</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-109.5,108,-109.5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-68.5,103,-25</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>103,-53.5,193,-53.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection>
<intersection>181 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>181,-60.5,181,-53.5</points>
<intersection>-60.5 13</intersection>
<intersection>-53.5 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>181,-60.5,200,-60.5</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>181 12</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-108.5,96,-76.5</points>
<intersection>-108.5 5</intersection>
<intersection>-87.5 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-87.5,98.5,-87.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96,-76.5,102,-76.5</points>
<intersection>96 0</intersection>
<intersection>102 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>102,-76.5,102,-74.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>96,-108.5,98.5,-108.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-122.5,88.5,-8</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-122.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-122.5,94.5,-122.5</points>
<intersection>88.5 0</intersection>
<intersection>94.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94.5,-127.5,94.5,-49</points>
<intersection>-127.5 9</intersection>
<intersection>-122.5 1</intersection>
<intersection>-110.5 7</intersection>
<intersection>-49 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>94.5,-49,200,-49</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>94.5 3</intersection>
<intersection>97.5 12</intersection>
<intersection>190.5 13</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>94.5,-110.5,98.5,-110.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>94.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>94.5,-127.5,101,-127.5</points>
<connection>
<GID>49</GID>
<name>IN_2</name></connection>
<intersection>94.5 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>97.5,-89.5,97.5,-49</points>
<intersection>-89.5 15</intersection>
<intersection>-49 5</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>190.5,-57,190.5,-49</points>
<intersection>-57 14</intersection>
<intersection>-49 5</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>190.5,-57,191.5,-57</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>190.5 13</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>97.5,-89.5,98.5,-89.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>97.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-93,107.5,-87.5</points>
<intersection>-93 2</intersection>
<intersection>-88.5 5</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-87.5,111,-87.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-93,107.5,-93</points>
<intersection>92.5 3</intersection>
<intersection>107.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>92.5,-102,92.5,-93</points>
<intersection>-102 7</intersection>
<intersection>-93 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>104.5,-88.5,107.5,-88.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>92.5,-102,98.5,-102</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>92.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-109,18.5,-106</points>
<intersection>-109 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-109,22.5,-109</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-106,18.5,-106</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-114.5,18,-111</points>
<intersection>-114.5 2</intersection>
<intersection>-111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-111,22.5,-111</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-114.5,18,-114.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-122.5,15.5,-22.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-122.5 9</intersection>
<intersection>-73.5 11</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>15.5,-122.5,184.5,-122.5</points>
<intersection>15.5 0</intersection>
<intersection>184.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>184.5,-122.5,184.5,-105.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-122.5 9</intersection>
<intersection>-112.5 14</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>13,-73.5,15.5,-73.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>184.5,-112.5,193.5,-112.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>184.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-113.5,7,-81.5</points>
<intersection>-113.5 5</intersection>
<intersection>-92.5 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-92.5,8.5,-92.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-81.5,12,-81.5</points>
<intersection>7 0</intersection>
<intersection>12 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>12,-81.5,12,-79.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>7,-113.5,8.5,-113.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-133.5,-1,-9</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-133.5,181.5,-133.5</points>
<intersection>-1 0</intersection>
<intersection>4.5 3</intersection>
<intersection>97.5 9</intersection>
<intersection>181.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4.5,-133.5,4.5,-94.5</points>
<intersection>-133.5 1</intersection>
<intersection>-115.5 7</intersection>
<intersection>-94.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4.5,-94.5,8.5,-94.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>4.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>4.5,-115.5,8.5,-115.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>4.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>181.5,-133.5,181.5,-101</points>
<intersection>-133.5 1</intersection>
<intersection>-109 12</intersection>
<intersection>-101 10</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>97.5,-133.5,97.5,-129.5</points>
<intersection>-133.5 1</intersection>
<intersection>-129.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>181.5,-101,193.5,-101</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>181.5 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>97.5,-129.5,101,-129.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>97.5 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>181.5,-109,185.5,-109</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>181.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-98,17.5,-92.5</points>
<intersection>-98 2</intersection>
<intersection>-93.5 5</intersection>
<intersection>-92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-92.5,21,-92.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-98,17.5,-98</points>
<intersection>8.5 3</intersection>
<intersection>17.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8.5,-107,8.5,-98</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>-98 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-93.5,17.5,-93.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-111.5,0.5,-101.5</points>
<intersection>-111.5 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-101.5,5,-101.5</points>
<intersection>-8 3</intersection>
<intersection>0.5 0</intersection>
<intersection>5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-111.5,0.5,-111.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>0.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-8,-101.5,-8,-73.5</points>
<intersection>-101.5 1</intersection>
<intersection>-100 7</intersection>
<intersection>-73.5 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>5,-105,5,-101.5</points>
<intersection>-105 5</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>5,-105,8.5,-105</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-8,-73.5,11,-73.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-8 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-8,-100,19.5,-100</points>
<intersection>-8 3</intersection>
<intersection>19.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>19.5,-100,19.5,-65.5</points>
<intersection>-100 7</intersection>
<intersection>-94.5 10</intersection>
<intersection>-65.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>19.5,-65.5,145.5,-65.5</points>
<intersection>19.5 8</intersection>
<intersection>57.5 13</intersection>
<intersection>101 12</intersection>
<intersection>145.5 15</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>19.5,-94.5,21,-94.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>19.5 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>101,-68.5,101,-65.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-65.5 9</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>57.5,-68.5,57.5,-65.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-65.5 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>145.5,-68,145.5,-65.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-65.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-93.5,28,-90</points>
<connection>
<GID>47</GID>
<name>N_in2</name></connection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-93.5,28,-93.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-88.5,118,-85</points>
<connection>
<GID>19</GID>
<name>N_in2</name></connection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,-88.5,118,-88.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-104,83.5,-96.5</points>
<intersection>-104 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-96.5,111,-96.5</points>
<intersection>83.5 0</intersection>
<intersection>98.5 4</intersection>
<intersection>111 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-104,83.5,-104</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>83.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,-96.5,111,-89.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>98.5,-100,98.5,-96.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-96.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-103.5,153,-100.5</points>
<intersection>-103.5 1</intersection>
<intersection>-100.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153,-103.5,157,-103.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149,-100.5,153,-100.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-109,152.5,-105.5</points>
<intersection>-109 2</intersection>
<intersection>-105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,-105.5,157,-105.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>152.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149,-109,152.5,-109</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>152.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-68,147.5,-22</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>147.5,-32.5,194,-32.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection>
<intersection>183 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>183,-37.5,183,-32.5</points>
<intersection>-37.5 19</intersection>
<intersection>-32.5 17</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>183,-37.5,203,-37.5</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>183 18</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-108,141.5,-76</points>
<intersection>-108 5</intersection>
<intersection>-87 1</intersection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-87,143,-87</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141.5,-76,146.5,-76</points>
<intersection>141.5 0</intersection>
<intersection>146.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>146.5,-76,146.5,-74</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>141.5,-108,143,-108</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-122,133.5,-5.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-122 1</intersection>
<intersection>-121.5 8</intersection>
<intersection>-27.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-122,139,-122</points>
<intersection>133.5 0</intersection>
<intersection>139 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>139,-122,139,-89</points>
<intersection>-122 1</intersection>
<intersection>-110 7</intersection>
<intersection>-89 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>139,-89,143,-89</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>139 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139,-110,143,-110</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>139 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>96.5,-121.5,133.5,-121.5</points>
<intersection>96.5 9</intersection>
<intersection>133.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>96.5,-126.5,96.5,-121.5</points>
<intersection>-126.5 10</intersection>
<intersection>-121.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>96.5,-126.5,101,-126.5</points>
<connection>
<GID>49</GID>
<name>IN_3</name></connection>
<intersection>96.5 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>133.5,-27.5,203,-27.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>133.5 0</intersection>
<intersection>192 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>192,-35.5,192,-27.5</points>
<intersection>-35.5 13</intersection>
<intersection>-27.5 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>192,-35.5,194,-35.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>192 12</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-92.5,152,-87</points>
<intersection>-92.5 2</intersection>
<intersection>-88 5</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,-87,155.5,-87</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>138,-92.5,152,-92.5</points>
<intersection>138 3</intersection>
<intersection>152 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>138,-101.5,138,-92.5</points>
<intersection>-101.5 7</intersection>
<intersection>-92.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>149,-88,152,-88</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>138,-101.5,143,-101.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>138 3</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-88,162.5,-84.5</points>
<connection>
<GID>28</GID>
<name>N_in2</name></connection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161.5,-88,162.5,-88</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>162.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-105,130.5,-95.5</points>
<intersection>-105 2</intersection>
<intersection>-95.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-95.5,155.5,-95.5</points>
<intersection>130.5 0</intersection>
<intersection>143 4</intersection>
<intersection>155.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118.5,-105,130.5,-105</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>130.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>155.5,-95.5,155.5,-89</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-95.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>143,-99.5,143,-95.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-95.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>163,-104.5,164.5,-104.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200.5,-32.5,200.5,-29.5</points>
<intersection>-32.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200.5,-29.5,203,-29.5</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>200.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-32.5,200.5,-32.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>200.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215.5,-28.5,215.5,-16.5</points>
<intersection>-28.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215.5,-16.5,258.5,-16.5</points>
<intersection>215.5 0</intersection>
<intersection>220 4</intersection>
<intersection>258.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,-28.5,215.5,-28.5</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>215.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>258.5,-21,258.5,-16.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>220,-24.5,220,-16.5</points>
<intersection>-24.5 5</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>220,-24.5,222.5,-24.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>220 4</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>198,-35.5,203,-35.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-46.5,219,-26.5</points>
<intersection>-46.5 3</intersection>
<intersection>-36.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-26.5,222.5,-26.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>209,-36.5,219,-36.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>219,-46.5,274,-46.5</points>
<intersection>219 0</intersection>
<intersection>274 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>274,-98,274,-46.5</points>
<intersection>-98 5</intersection>
<intersection>-46.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>274,-98,278.5,-98</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>274 4</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-24.5,238,-24.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>228.5 7</intersection>
<intersection>236 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>236,-96,236,-24.5</points>
<intersection>-96 9</intersection>
<intersection>-65 6</intersection>
<intersection>-37 4</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>236,-37,239.5,-37</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>236 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>236,-65,250.5,-65</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>236 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>228.5,-25.5,228.5,-24.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>236,-96,259.5,-96</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>236 3</intersection>
<intersection>236.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>236.5,-153.5,236.5,-96</points>
<intersection>-153.5 13</intersection>
<intersection>-115.5 11</intersection>
<intersection>-96 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>236.5,-115.5,253.5,-115.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>236.5 10</intersection>
<intersection>246 14</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>236.5,-153.5,254.5,-153.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>236.5 10</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>246,-122,246,-115.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-115.5 11</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-53.5,197.5,-51</points>
<intersection>-53.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197.5,-51,200,-51</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-53.5,197.5,-53.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>197.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-58.5,197.5,-57</points>
<intersection>-58.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197.5,-58.5,200,-58.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>197.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195.5,-57,197.5,-57</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>197.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>206,-50,231.5,-50</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>214 5</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>231.5,-50,231.5,-26.5</points>
<intersection>-50 1</intersection>
<intersection>-26.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>231.5,-26.5,238,-26.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>214,-53,214,-50</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-50 1</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-98,208,-55</points>
<intersection>-98 3</intersection>
<intersection>-59.5 2</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208,-55,214,-55</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>206,-59.5,208,-59.5</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>208,-98,259.5,-98</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-117,229.5,-39</points>
<intersection>-117 5</intersection>
<intersection>-67 3</intersection>
<intersection>-54 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>229.5,-39,239.5,-39</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-54,229.5,-54</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>229.5,-67,250.5,-67</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>229.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>229.5,-117,253.5,-117</points>
<intersection>229.5 0</intersection>
<intersection>230 6</intersection>
<intersection>240.5 8</intersection>
<intersection>253.5 9</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>230,-155.5,230,-117</points>
<intersection>-155.5 7</intersection>
<intersection>-117 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>230,-155.5,254.5,-155.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>230 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>240.5,-124,240.5,-117</points>
<intersection>-124 10</intersection>
<intersection>-117 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>253.5,-117.5,253.5,-117</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>-117 5</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>240.5,-124,246,-124</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>240.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-80,192,-74.5</points>
<intersection>-80 2</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-74.5,194,-74.5</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190,-80,192,-80</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>192 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,-86.5,192.5,-85</points>
<intersection>-86.5 1</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192.5,-86.5,194.5,-86.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>192.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>190.5,-85,192.5,-85</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-73.5,239.5,-73.5</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>209 4</intersection>
<intersection>239.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>239.5,-73.5,239.5,-41</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>209,-75.5,209,-73.5</points>
<intersection>-75.5 5</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>209,-75.5,210,-75.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>209 4</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>202,-119.5,202,-77.5</points>
<intersection>-119.5 3</intersection>
<intersection>-87.5 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202,-77.5,210,-77.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>202 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-87.5,202,-87.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>202 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>202,-119.5,253.5,-119.5</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>202 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225.5,-157.5,225.5,-69</points>
<intersection>-157.5 3</intersection>
<intersection>-126 4</intersection>
<intersection>-76.5 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225.5,-69,250.5,-69</points>
<connection>
<GID>86</GID>
<name>IN_2</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>216,-76.5,225.5,-76.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>225.5,-157.5,254.5,-157.5</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>225.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>225.5,-126,246,-126</points>
<connection>
<GID>98</GID>
<name>IN_2</name></connection>
<intersection>225.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-105.5,191,-103</points>
<intersection>-105.5 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-103,193.5,-103</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>191 0</intersection>
<intersection>192.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,-105.5,191,-105.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>191 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>192.5,-128,192.5,-103</points>
<intersection>-128 4</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>192.5,-128,246,-128</points>
<connection>
<GID>98</GID>
<name>IN_3</name></connection>
<intersection>192.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-110.5,191.5,-109</points>
<intersection>-110.5 1</intersection>
<intersection>-109 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-110.5,193.5,-110.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>189.5,-109,191.5,-109</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>199.5,-102,250.5,-102</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>208.5 4</intersection>
<intersection>250.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>250.5,-102,250.5,-71</points>
<connection>
<GID>86</GID>
<name>IN_3</name></connection>
<intersection>-102 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>208.5,-106,208.5,-102</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>-102 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204,-111.5,204,-108</points>
<intersection>-111.5 2</intersection>
<intersection>-108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204,-108,208.5,-108</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>204 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>199.5,-111.5,204,-111.5</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>204 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-159.5,218.5,-107</points>
<intersection>-159.5 1</intersection>
<intersection>-107 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-159.5,254.5,-159.5</points>
<connection>
<GID>96</GID>
<name>IN_3</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214.5,-107,218.5,-107</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-117.5,269,-104</points>
<intersection>-117.5 2</intersection>
<intersection>-104 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269,-104,278.5,-104</points>
<connection>
<GID>97</GID>
<name>IN_3</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>259.5,-117.5,269,-117.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,-102,272,-97</points>
<intersection>-102 1</intersection>
<intersection>-97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272,-102,278.5,-102</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<intersection>272 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265.5,-97,272,-97</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>272 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,-100,247,-23</points>
<intersection>-100 3</intersection>
<intersection>-25.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,-23,258.5,-23</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,-25.5,247,-25.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>247,-100,278.5,-100</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252,-39,252,-25</points>
<intersection>-39 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252,-25,258.5,-25</points>
<connection>
<GID>71</GID>
<name>IN_2</name></connection>
<intersection>252 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>245.5,-39,252,-39</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>252 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257.5,-68,257.5,-27</points>
<intersection>-68 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257.5,-27,258.5,-27</points>
<connection>
<GID>71</GID>
<name>IN_3</name></connection>
<intersection>257.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>256.5,-68,257.5,-68</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>257.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-24,269,-23.5</points>
<intersection>-24 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269,-23.5,273,-23.5</points>
<connection>
<GID>99</GID>
<name>N_in1</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>265.5,-24,269,-24</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-101,287,-100.5</points>
<intersection>-101 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>287,-100.5,289,-100.5</points>
<connection>
<GID>100</GID>
<name>N_in0</name></connection>
<intersection>287 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>285.5,-101,287,-101</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>287 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>260.5,-156.5,267.5,-156.5</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<connection>
<GID>101</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 1>
<page 2>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 2>
<page 3>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 3>
<page 4>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 4>
<page 5>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 5>
<page 6>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 6>
<page 7>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 7>
<page 8>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 8>
<page 9>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 9></circuit>