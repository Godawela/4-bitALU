<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-14.4194,17.0221,171.056,-76.3808</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>20,-13</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>21,-19</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>21,-36</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_XOR2</type>
<position>38.5,-14</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>39,-25</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>54,-17.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_OR2</type>
<position>68.5,-24</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>80,-23.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AI_XOR2</type>
<position>66,-7</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>77,-7</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-13,35.5,-13</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>33.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-24,33.5,-13</points>
<intersection>-24 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33.5,-24,36,-24</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>33.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-26,29,-15</points>
<intersection>-26 3</intersection>
<intersection>-19 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-19,29,-19</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-15,35.5,-15</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-26,36,-26</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-14,60,-14</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>51 4</intersection>
<intersection>60 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60,-14,60,-8</points>
<intersection>-14 1</intersection>
<intersection>-8 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>51,-16.5,51,-14</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>60,-8,63,-8</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>60 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-36,49,-18.5</points>
<intersection>-36 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-18.5,51,-18.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>46 3</intersection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-36,49,-36</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46,-18.5,46,-6</points>
<intersection>-18.5 1</intersection>
<intersection>-6 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46,-6,63,-6</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>46 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-23,60.5,-17.5</points>
<intersection>-23 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-23,65.5,-23</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-17.5,60.5,-17.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-25,65.5,-25</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-24,79,-24</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>79 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>79,-24,79,-23.5</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-7,76,-7</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 1>
<page 2>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 2>
<page 3>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 3>
<page 4>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 4>
<page 5>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 5>
<page 6>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 6>
<page 7>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 7>
<page 8>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 8>
<page 9>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 9></circuit>