<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-5.94999,33.5692,240.831,-90.7063</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>69,-6.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>12.5,-47</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>80,-24</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>80,-36.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>80,-45</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>80.5,-7</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>81.5,2</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AI_XOR2</type>
<position>94.5,-23.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AE_OR2</type>
<position>88,-39.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>98.5,-19</position>
<input>
<ID>N_in0</ID>10 </input>
<input>
<ID>N_in1</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>112.5,-6.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AI_XOR2</type>
<position>123.5,-24</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AI_XOR2</type>
<position>136,-24</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>123.5,-36.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND2</type>
<position>123.5,-45</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR2</type>
<position>137.5,-40.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR2</type>
<position>124,-7</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>125,2</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>140,-19.5</position>
<input>
<ID>N_in1</ID>40 </input>
<input>
<ID>N_in2</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>157,-6</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>168,-23.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AI_XOR2</type>
<position>180.5,-23.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>168,-36</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>168,-44.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_OR2</type>
<position>182,-40</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AI_XOR2</type>
<position>168.5,-6.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>169.5,2.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>184.5,-19</position>
<input>
<ID>N_in1</ID>41 </input>
<input>
<ID>N_in2</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>198,-31.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>41 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>187.5,-40</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>192.5,0</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>1 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>30 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>196.5,1.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>22.5,-11.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AI_XOR2</type>
<position>33.5,-29</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>201.5,-36.5</position>
<gparam>LABEL_TEXT Output</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AI_XOR2</type>
<position>46,-29</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>33.5,-41.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>187.5,-43</position>
<gparam>LABEL_TEXT C3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>33.5,-50</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>140.5,-44</position>
<gparam>LABEL_TEXT C2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AE_OR2</type>
<position>47.5,-45.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>91.5,-43</position>
<gparam>LABEL_TEXT C1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AI_XOR2</type>
<position>34,-12</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>51.5,-48</position>
<gparam>LABEL_TEXT C0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>35,-3</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>19,-11.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>50,-24.5</position>
<input>
<ID>N_in1</ID>38 </input>
<input>
<ID>N_in2</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>30.5,-3</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>123.5,-62</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>32 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>64.5,-6.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>77.5,2.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>108,-6.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>120.5,2</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>153,-5.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>165.5,3</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>9,-46.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>10,-50</position>
<gparam>LABEL_TEXT Add 0 / Sub 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>50,-21.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>98,-16.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>137.5,-19</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>184,-16.5</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-4,84.5,6.5</points>
<intersection>-4 7</intersection>
<intersection>0 6</intersection>
<intersection>6.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>84.5,6.5,186.5,6.5</points>
<intersection>84.5 0</intersection>
<intersection>186.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>186.5,0,186.5,6.5</points>
<intersection>0 5</intersection>
<intersection>6.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>186.5,0,189.5,0</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>186.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>81.5,0,84.5,0</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>81.5,-4,84.5,-4</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-44,75.5,-12</points>
<intersection>-44 5</intersection>
<intersection>-23 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-23,77,-23</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-12,80.5,-12</points>
<intersection>75.5 0</intersection>
<intersection>80.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80.5,-12,80.5,-10</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>75.5,-44,77,-44</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-58,67.5,-12</points>
<intersection>-58 1</intersection>
<intersection>-12 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-58,104.5,-58</points>
<intersection>67.5 0</intersection>
<intersection>73 3</intersection>
<intersection>77 9</intersection>
<intersection>104.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73,-58,73,-25</points>
<intersection>-58 1</intersection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>67.5,-12,69,-12</points>
<intersection>67.5 0</intersection>
<intersection>69 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>73,-25,77,-25</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>73 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>69,-12,69,-8.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-12 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>104.5,-62,104.5,-58</points>
<intersection>-62 10</intersection>
<intersection>-58 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>77,-58,77,-46</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>104.5,-62,120.5,-62</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>104.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-28.5,86,-22.5</points>
<intersection>-28.5 2</intersection>
<intersection>-24 5</intersection>
<intersection>-22.5 8</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-28.5,86,-28.5</points>
<intersection>70.5 3</intersection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-37.5,70.5,-28.5</points>
<intersection>-37.5 7</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>83,-24,86,-24</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>70.5,-37.5,77,-37.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>70.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>86,-22.5,91.5,-22.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-45.5,63.5,-32</points>
<intersection>-45.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-32,91.5,-32</points>
<intersection>63.5 0</intersection>
<intersection>74 4</intersection>
<intersection>91.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-45.5,63.5,-45.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91.5,-32,91.5,-24.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>74,-35.5,74,-32</points>
<intersection>-35.5 5</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>74,-35.5,77,-35.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>74 4</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-38.5,84,-36.5</points>
<intersection>-38.5 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-38.5,85,-38.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-36.5,84,-36.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-45,84,-40.5</points>
<intersection>-45 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-40.5,85,-40.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-45,84,-45</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-23.5,98,-19</points>
<intersection>-23.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,-19,98,-19</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-23.5,98,-23.5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-39.5,130.5,-36.5</points>
<intersection>-39.5 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-39.5,134.5,-39.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>130.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126.5,-36.5,130.5,-36.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-45,130,-41.5</points>
<intersection>-45 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-41.5,134.5,-41.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126.5,-45,130,-45</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-4,130,10.5</points>
<intersection>-4 7</intersection>
<intersection>0 6</intersection>
<intersection>10.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>130,10.5,184.5,10.5</points>
<intersection>130 0</intersection>
<intersection>184.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>184.5,1,184.5,10.5</points>
<intersection>1 5</intersection>
<intersection>10.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>184.5,1,189.5,1</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>184.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>125,0,130,0</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>125,-4,130,-4</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-44,119,-12</points>
<intersection>-44 5</intersection>
<intersection>-23 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-23,120.5,-23</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,-12,124,-12</points>
<intersection>119 0</intersection>
<intersection>124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124,-12,124,-10</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>119,-44,120.5,-44</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-58,111,-12</points>
<intersection>-58 1</intersection>
<intersection>-12 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-58,116.5,-58</points>
<intersection>111 0</intersection>
<intersection>116.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116.5,-61,116.5,-25</points>
<intersection>-61 9</intersection>
<intersection>-58 1</intersection>
<intersection>-46 7</intersection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>111,-12,112.5,-12</points>
<intersection>111 0</intersection>
<intersection>112.5 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>116.5,-25,120.5,-25</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>116.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>112.5,-12,112.5,-8.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-12 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>116.5,-46,120.5,-46</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>116.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>116.5,-61,120.5,-61</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<intersection>116.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-28.5,129.5,-23</points>
<intersection>-28.5 2</intersection>
<intersection>-24 5</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-23,133,-23</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-28.5,129.5,-28.5</points>
<intersection>114.5 3</intersection>
<intersection>129.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114.5,-37.5,114.5,-28.5</points>
<intersection>-37.5 7</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>126.5,-24,129.5,-24</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114.5,-37.5,120.5,-37.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>114.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-44.5,40.5,-41.5</points>
<intersection>-44.5 1</intersection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-44.5,44.5,-44.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-41.5,40.5,-41.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-50,40,-46.5</points>
<intersection>-50 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-46.5,44.5,-46.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-50,40,-50</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-9,35,5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,5,188,5</points>
<intersection>35 0</intersection>
<intersection>188 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>188,-1,188,5</points>
<intersection>-1 3</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>188,-1,189.5,-1</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>188 2</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-49,29,-17</points>
<intersection>-49 5</intersection>
<intersection>-28 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-28,30.5,-28</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-17,34,-17</points>
<intersection>29 0</intersection>
<intersection>34 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-17,34,-15</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>29,-49,30.5,-49</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-63,21,-17</points>
<intersection>-63 1</intersection>
<intersection>-17 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-63,120.5,-63</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection>
<intersection>26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-63,26.5,-30</points>
<intersection>-63 1</intersection>
<intersection>-51 7</intersection>
<intersection>-30 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21,-17,22.5,-17</points>
<intersection>21 0</intersection>
<intersection>22.5 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-30,30.5,-30</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>26.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>22.5,-17,22.5,-13.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-17 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>26.5,-51,30.5,-51</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>26.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-33.5,39.5,-28</points>
<intersection>-33.5 2</intersection>
<intersection>-29 5</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-28,43,-28</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-33.5,39.5,-33.5</points>
<intersection>30.5 3</intersection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-42.5,30.5,-33.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>36.5,-29,39.5,-29</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-47,22.5,-37</points>
<intersection>-47 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-37,27,-37</points>
<intersection>14 3</intersection>
<intersection>22.5 0</intersection>
<intersection>27 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-47,22.5,-47</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-37,14,-9</points>
<intersection>-37 1</intersection>
<intersection>-35.5 7</intersection>
<intersection>-9 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>27,-40.5,27,-37</points>
<intersection>-40.5 5</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>27,-40.5,30.5,-40.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>27 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>14,-9,33,-9</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>14 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>14,-35.5,41.5,-35.5</points>
<intersection>14 3</intersection>
<intersection>41.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>41.5,-35.5,41.5,-1</points>
<intersection>-35.5 7</intersection>
<intersection>-30 10</intersection>
<intersection>-1 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>41.5,-1,167.5,-1</points>
<intersection>41.5 8</intersection>
<intersection>79.5 13</intersection>
<intersection>123 12</intersection>
<intersection>167.5 15</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>41.5,-30,43,-30</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>41.5 8</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>123,-4,123,-1</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-1 9</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>79.5,-4,79.5,-1</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-1 9</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>167.5,-3.5,167.5,-1</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>-1 9</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-29,50,-25.5</points>
<connection>
<GID>58</GID>
<name>N_in2</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-29,50,-29</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-24,140,-20.5</points>
<connection>
<GID>23</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,-24,140,-24</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-39.5,105.5,-32</points>
<intersection>-39.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-32,133,-32</points>
<intersection>105.5 0</intersection>
<intersection>120.5 4</intersection>
<intersection>133 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-39.5,105.5,-39.5</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>105.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>133,-32,133,-25</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>120.5,-35.5,120.5,-32</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-32 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-39,175,-36</points>
<intersection>-39 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-39,179,-39</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171,-36,175,-36</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-44.5,174.5,-41</points>
<intersection>-44.5 2</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174.5,-41,179,-41</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>174.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171,-44.5,174.5,-44.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>174.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-3.5,169.5,8</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>8 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>169.5,8,183.5,8</points>
<intersection>169.5 0</intersection>
<intersection>183.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>183.5,2,183.5,8</points>
<intersection>2 11</intersection>
<intersection>8 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>183.5,2,189.5,2</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>183.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-43.5,163.5,-11.5</points>
<intersection>-43.5 5</intersection>
<intersection>-22.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-22.5,165,-22.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-11.5,168.5,-11.5</points>
<intersection>163.5 0</intersection>
<intersection>168.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>168.5,-11.5,168.5,-9.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>163.5,-43.5,165,-43.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-57.5,155.5,-11.5</points>
<intersection>-57.5 1</intersection>
<intersection>-57 8</intersection>
<intersection>-11.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,-57.5,161,-57.5</points>
<intersection>155.5 0</intersection>
<intersection>161 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>161,-57.5,161,-24.5</points>
<intersection>-57.5 1</intersection>
<intersection>-45.5 7</intersection>
<intersection>-24.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>155.5,-11.5,157,-11.5</points>
<intersection>155.5 0</intersection>
<intersection>157 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>161,-24.5,165,-24.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>161 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>157,-11.5,157,-8</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>161,-45.5,165,-45.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>161 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118.5,-57,155.5,-57</points>
<intersection>118.5 9</intersection>
<intersection>155.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>118.5,-60,118.5,-57</points>
<intersection>-60 10</intersection>
<intersection>-57 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>118.5,-60,120.5,-60</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<intersection>118.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-28,174,-22.5</points>
<intersection>-28 2</intersection>
<intersection>-23.5 5</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,-22.5,177.5,-22.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-28,174,-28</points>
<intersection>160 3</intersection>
<intersection>174 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>160,-37,160,-28</points>
<intersection>-37 7</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>171,-23.5,174,-23.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>160,-37,165,-37</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>160 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-23.5,184.5,-20</points>
<connection>
<GID>33</GID>
<name>N_in2</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183.5,-23.5,184.5,-23.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-40.5,152.5,-31</points>
<intersection>-40.5 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,-31,177.5,-31</points>
<intersection>152.5 0</intersection>
<intersection>165 4</intersection>
<intersection>177.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-40.5,152.5,-40.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>152.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>177.5,-31,177.5,-24.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-31 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>165,-35,165,-31</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,-40,186.5,-40</points>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-32.5,113.5,-27</points>
<intersection>-32.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113.5,-32.5,195,-32.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-27,113.5,-27</points>
<intersection>52.5 3</intersection>
<intersection>113.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-27,52.5,-24.5</points>
<intersection>-27 2</intersection>
<intersection>-24.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51,-24.5,52.5,-24.5</points>
<connection>
<GID>58</GID>
<name>N_in1</name></connection>
<intersection>52.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-31.5,147,-16.5</points>
<intersection>-31.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-31.5,195,-31.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>101,-16.5,147,-16.5</points>
<intersection>101 3</intersection>
<intersection>147 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101,-19,101,-16.5</points>
<intersection>-19 4</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>99.5,-19,101,-19</points>
<connection>
<GID>13</GID>
<name>N_in1</name></connection>
<intersection>101 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158,-30.5,158,-19.5</points>
<intersection>-30.5 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,-30.5,195,-30.5</points>
<connection>
<GID>35</GID>
<name>IN_2</name></connection>
<intersection>158 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-19.5,158,-19.5</points>
<connection>
<GID>23</GID>
<name>N_in1</name></connection>
<intersection>158 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-29.5,190,-19</points>
<intersection>-29.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-29.5,195,-29.5</points>
<connection>
<GID>35</GID>
<name>IN_3</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185.5,-19,190,-19</points>
<connection>
<GID>33</GID>
<name>N_in1</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 1>
<page 2>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 2>
<page 3>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 3>
<page 4>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 4>
<page 5>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 5>
<page 6>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 6>
<page 7>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 7>
<page 8>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 8>
<page 9>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 9></circuit>