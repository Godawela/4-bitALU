<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>5.05692,20.3307,83.4694,-61.6299</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>18,-10</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>19,-18.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>19,-25.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>19,-33</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,-10</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>27,-18.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_SMALL_INVERTER</type>
<position>27.5,-25.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_SMALL_INVERTER</type>
<position>27.5,-33</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>39.5,-9</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>39,-17.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>38,-27.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AI_XOR2</type>
<position>53.5,-33.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>53.5,-24</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AI_XOR2</type>
<position>53,-14.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AI_XOR2</type>
<position>52.5,-6</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>67.5,-33.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>67.5,-23.5</position>
<input>
<ID>N_in2</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>67.5,-14.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>67,-6</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>EE_VDD</type>
<position>26.5,-1.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>12.5,-10</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>12,-18</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>12,-24.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>12,-32.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-10,24,-10</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-18.5,25,-18.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-25.5,25.5,-25.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-33,25.5,-33</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-33.5,66.5,-33.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-24.5,67.5,-24</points>
<connection>
<GID>34</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-24,67.5,-24</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-14.5,66.5,-14.5</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<connection>
<GID>28</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-6,66,-6</points>
<connection>
<GID>38</GID>
<name>N_in0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-34.5,40,-33</points>
<intersection>-34.5 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-34.5,50.5,-34.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-33,40,-33</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-31.5,33,-25.5</points>
<intersection>-31.5 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-31.5,50.5,-31.5</points>
<intersection>33 0</intersection>
<intersection>35 4</intersection>
<intersection>50.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-25.5,33,-25.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-31.5,50.5,-25</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>35,-31.5,35,-28.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-32.5,43.5,-27.5</points>
<intersection>-32.5 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-32.5,50.5,-32.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-27.5,43.5,-27.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-22.5,48,-22.5</points>
<intersection>33.5 5</intersection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48,-22.5,48,-15.5</points>
<intersection>-22.5 1</intersection>
<intersection>-15.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48,-15.5,50,-15.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>33.5,-22.5,33.5,-18.5</points>
<intersection>-22.5 1</intersection>
<intersection>-18.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>29,-18.5,36,-18.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>33.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-24,44,-17.5</points>
<intersection>-24 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-24,44,-24</points>
<intersection>35 4</intersection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-17.5,50.5,-17.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>44 0</intersection>
<intersection>50.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-23,50.5,-17.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-17.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>35,-26.5,35,-24</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-13.5,46,-9</points>
<intersection>-13.5 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-13.5,50,-13.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-9,46,-9</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>44 3</intersection>
<intersection>46 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-14,44,-9</points>
<intersection>-14 4</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-14,44,-14</points>
<intersection>36 5</intersection>
<intersection>44 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>36,-16.5,36,-14</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-14 4</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-12.5,34.5,-10</points>
<intersection>-12.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-12.5,49.5,-12.5</points>
<intersection>34.5 0</intersection>
<intersection>49.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-10,36.5,-10</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-12.5,49.5,-7</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-3.5,26.5,-2.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-3.5,45,-3.5</points>
<intersection>26.5 0</intersection>
<intersection>36.5 3</intersection>
<intersection>45 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>45,-5,45,-3.5</points>
<intersection>-5 4</intersection>
<intersection>-3.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>36.5,-8,36.5,-3.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45,-5,49.5,-5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>45 2</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 1>
<page 2>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 2>
<page 3>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 3>
<page 4>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 4>
<page 5>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 5>
<page 6>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 6>
<page 7>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 7>
<page 8>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 8>
<page 9>
<PageViewport>0,37.7538,139.4,-107.954</PageViewport></page 9></circuit>